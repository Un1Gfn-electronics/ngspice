.title voltage divider netlist
.options TEMP=27 TNOM=27

V1 in  0   1
R1 out in  1k
R2 0   out 2k

.tran 1ns 3ns

.end
