* https://www.youtube.com/watch?v=_vKeaPHXF9U&list=PLBlnK6fEyqRiw-GZRqfnlVIBz9dxrqHJS&index=15

.title V-I Characteristics of PN Junction Diode

V1 a 0 dc 0 PULSE( 0v 1v 0s 100s )

D1 a 0 Silicon area=1.0 
* .model Silicon D( IS=100uA RS=333 BV=100V VJ=100v PHP=100v )
.model Silicon D( IS=100uA EG=1.11 BV=0.1V VJ=0.2v PHP=0.3v )
.save all @d1[id]

.tran 10ms 100s

.control
  run
  plot @d1[id] vs a
  * plot @d1[id] vs a xlimit -250mV 0 ylimit -110mA 0
.endc

.end
