* https://www.youtube.com/watch?v=_vKeaPHXF9U&list=PLBlnK6fEyqRiw-GZRqfnlVIBz9dxrqHJS&index=15

.title V-I Characteristics of PN Junction Diode

V1   a 0 dc 0 PULSE( 0v 1v 0s 1s )

.model Silicon D(EG=1.11)
D_Si a 0 Silicon area=1.0

* id is current_of_diode
.save all @D_Si[id]

.tran 10us 1s

.control
  run
  plot @D_Si[id] vs a nointerp
  plot @D_Si[id] vs a ylimit 0 100uA nointerp
.endc

.end
