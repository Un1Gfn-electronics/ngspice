* https://wiki.analog.com/university/courses/electronics/electronics-lab-27
* ngspice -nb inv.cir
.title TTL Inverter

.include 2N3904.SP3
.include SSM2212.cir
.include 1N914.mod

* Input current steering stage
.SUBCKT ICSS   Vcc Vin             Q1C
  R1 Vcc o       100k
  Q1 Q1C o Vin 2N3904
.ENDS

* Phase splitting stage
.SUBCKT PSS    Vcc GND Vin         Vo1 Vo2
  R2 Vcc Vo1     2200
  R3 GND Vo2     470
  Q2 Vo1 Vin Vo2 2N3904
.ENDS

* Output Stage
.SUBCKT OS     Vcc GND Vi1 Vi2     Vout
  *
  R4   Vcc Q4C                      100
  D1   Q4E Vout                     FDLL914B
  *
  *    Q4C Q4B Q4E   Q3E Q3B Q3C
  Xssm Q4C Vi1 Q4E   GND Vi2 Vout   SSM2212
  *
.ENDS

Vx   x 0 0v
VC Vcc 0 6v

XUicss         Vcc x             Q1C       ICSS
XUpss          Vcc 0 Q1C         Vo1 Vo2   PSS
XUos           Vcc 0 Vo1 Vo2     y         OS

.control
  foreach xx 0 6v
    alter Vx=$xx
    op
    echo
    echo
    echo
    print x y
    echo
    echo
    echo
    shell read -r
  end
.endc

.end
