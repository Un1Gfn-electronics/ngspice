* https://wiki.analog.com/university/courses/electronics/electronics-lab-27
* ngspice -nb inv.cir
.title TTL Inverter

.include 2N3904.SP3

* Input current steering stage
.SUBCKT ICSS   Vcc Vin             Q1C
  R1 Vcc o       100k
  Q1 Q1C o Vin 2N3904
.ENDS


* Phase splitting stage
.SUBCKT PSS    Vcc GND Vin         Vo1 Vo2
.ENDS

* Output Stage
.SUBCKT OS     Vcc GND Vi1 Vi2     Vout 
.ENDS

Vx   x 0 0v
VC Vcc 0 6v
VG GND 0 0v

XUicss         Vcc x               Q1C       ICSS
XUpss          Vcc GND Q1C         Vo1 Vo2   PSS
XUos           Vcc GND Vo1 Vo2     y         OS

.control
  foreach xx 0 6v
      alter Vx=$xx
      * op
      echo
      echo
      echo
      * print x y
      echo
      echo
      echo
      shell read -r
    end
  end
.endc