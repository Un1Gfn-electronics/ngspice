* https://wiki.analog.com/university/courses/electronics/electronics-lab-27
* ngspice -nb inv.cir
.title TTL Inverter
.options TEMP=27 TNOM=27 WARN=1

.include 2N3904.SP3
.include SSM2212.cir
.include 1N914.mod

* https://sourceforge.net/p/ngspice/discussion/133842/thread/80d38e4d/#897d
.param   HIGH=6v
.csparam HIGH={HIGH}

* Input current steering stage
.SUBCKT ICSS   Vcc Vin             Q1C
  R1 Vcc o       100k
  Q1 Q1C o Vin 2N3904
.ENDS

* Phase splitting stage
.SUBCKT PSS    Vcc GND Vin         Vo1 Vo2
  R2 Vcc Vo1     2200
  R3 GND Vo2     470
  Q2 Vo1 Vin Vo2 2N3904
.ENDS

* Output Stage
.SUBCKT OS     Vcc GND Vi1 Vi2     Vout
  *
  R4   Vcc Q4C                      100
  D1   Q4E Vout                     FDLL914B
  *
  *    Q4C Q4B Q4E   Q3E Q3B Q3C
  Xssm Q4C Vi1 Q4E   GND Vi2 Vout   SSM2212
  *
.ENDS

* Vx   x 0 0v dc 0 PWL(0s 0v 1e-8s {HIGH})
Vx   x 0 0v dc 0 PULSE(0v {HIGH} 0 1e-8 1e-8 200e-8 402e-8)
VC Vcc 0 {HIGH}

XUicss         Vcc x             Q1C       ICSS
XUpss          Vcc 0 Q1C         Vo1 Vo2   PSS
XUos           Vcc 0 Vo1 Vo2     y         OS

.control
  tran 0.1e-8 803e-8
  print x[length(x)-1] y[length(y)-1]
  * plot x y pointplot
  * plot x y
  let shift={HIGH*1.01}
  plot x-shift y
  * plot x
  * plot y
.endc

.end
