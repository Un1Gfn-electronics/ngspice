.title Load Line Analysis (Numerical Problem)
.options TEMP=27 TNOM=27

V1 a 0 10v
R1 a b 1kOhm

B1 b 0 I=v(b)/v(c)
Vx c 0 dc 0

.save all @R1[i]

.dc Vx 1v 1e5v 1v

.control
  run
  plot @R1[i] vs b nointerp ylimit 0mA 11mA xlimit 0v 15v
.endc

.end
