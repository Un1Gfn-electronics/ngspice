.title Load Line Analysis (Numerical Problem)
.options TEMP=27 TNOM=27

V1 a 0 10v
R1 a b 1kOhm
B1 b 0 I=v(b)/v(c)
Vx c 0 dc 1e5v

V2   m 0 dc 0v
D_Si m 0 Silicon area=1.0
.model Silicon D(EG=1.11 BV=40)

.save all
.save @R1[i]
.save @D_Si[id]

.control
  *
  dc Vx   1v  1e5v  100v
  dc V2   0v    1v   10mV
  *
  dc Vx   1v  111v  100mv
  dc V2 710mV 720mV 100uV
  *
  * plot dc1.@R1[i]    vs dc1.b ylimit 0mA 11mA xlimit 0v 15v pointplot nointerp
  * plot dc2.@D_Si[id] vs dc2.m ylimit 0mA 11mA xlimit 0v 15v pointplot nointerp
  plot dc1.@R1[i] vs dc1.b dc2.@D_Si[id] vs dc2.m ylimit 0mA 11mA xlimit   0v   15v  pointplot nointerp
  plot dc3.@R1[i] vs dc3.b dc4.@D_Si[id] vs dc4.m ylimit 9mA 10mA xlimit 700mV 800mV pointplot nointerp
.endc

.end
