* https://wiki.analog.com/university/courses/electronics/electronics-lab-27
* ngspice -nb inv.cir
.title TTL Inverter
.options TEMP=27 TNOM=27 WARN=1

.include 2N3904.SP3
.include SSM2212.cir
.include 1N914.mod

* https://sourceforge.net/p/ngspice/discussion/133842/thread/80d38e4d/#897d
.param   HIGH=6v
.csparam HIGH={HIGH}

* Input current steering stage
.SUBCKT ICSS   Vcc Vin             Q1C
  R1 Vcc o       100k
  Q1 Q1C o Vin 2N3904
.ENDS

* Phase splitting stage
.SUBCKT PSS    Vcc GND Vin         Vo1 Vo2
  R2 Vcc Vo1     2200
  R3 GND Vo2     470
  Q2 Vo1 Vin Vo2 2N3904
.ENDS

* Output Stage
.SUBCKT OS     Vcc GND Vi1 Vi2     Vout
  *
  R4   Vcc Q4C                      100
  D1   Q4E Vout                     FDLL914B
  *
  *    Q4C Q4B Q4E   Q3E Q3B Q3C
  Xssm Q4C Vi1 Q4E   GND Vi2 Vout   SSM2212
  *
.ENDS

* Vx   x 0 0v dc 0 PWL(0s 0v 1e-8s {HIGH})
Vx   x 0 0v dc 0 PULSE(0v {HIGH} 0 1e-8 1e-8 200e-8 402e-8)
V0 Vcc 0 {HIGH}

.SUBCKT INV   Vcc GND x         y
  XUicss      Vcc x             Q1C       ICSS
  XUpss       Vcc GND Q1C       Vo1 Vo2   PSS
  XUos        Vcc GND Vo1 Vo2   y         OS
.ENDS

XNAND1   Vcc GND x  y1   INV
XNAND2   Vcc GND y1 y2   INV
XNAND3   Vcc GND y2 y3   INV
XNAND4   Vcc GND y3 y4   INV
XNAND5   Vcc GND y4 y5   INV
XNAND6   Vcc GND y5 y6   INV
XNAND7   Vcc GND y6 y7   INV
XNAND8   Vcc GND y7 y8   INV

.control

  tran 0.1e-8 1000e-8

  * plot x
  * plot y
  * plot x y
  * plot x y pointplot

  * print x[length(x)-1] y[length(y)-1]

  * let shift={HIGH*1.01}
  * plot x-shift y

  plot
  + x
  + y1+0.1*0.5
  + y2+0.2*0.5
  + y3+0.3*0.5
  + y4+0.4*0.5
  + y5+0.5*0.5
  + y6+0.6*0.5
  + y7+0.7*0.5
  + y8+0.8*0.5

.endc

.end
