* https://www.youtube.com/watch?v=_vKeaPHXF9U&list=PLBlnK6fEyqRiw-GZRqfnlVIBz9dxrqHJS&index=15

.title V-I Characteristics of PN Junction Diode

V1   a 0 dc 0 PULSE( 0v 1v 0s 100s )

.model Silicon   D(EG=1.11)
.model 1N34A D(bv=75 cjo=0.5e-12 eg=0.67 ibv=18e-3 is=2e-7 rs=7 n=1.3 vj=0.1 m=0.27)

D_Si a 0 Silicon   area=1.0
D_Ge a 0 1N34A area=1.0

.save all
.save @D_Si[id]
.save @D_Ge[id]

.tran 10ms 100s

.control
  run
  plot @D_Si[id] vs a
  plot @D_Ge[id] vs a
  * plot @D_Si[id] @D_Ge[id] vs a
  * plot @d1[id] vs a xlimit -2V 0 ylimit -110mA 0
.endc

.end
