* https://www.youtube.com/watch?v=_vKeaPHXF9U&list=PLBlnK6fEyqRiw-GZRqfnlVIBz9dxrqHJS&index=15

.title V-I Characteristics of PN Junction Diode

V1 a 0 dc 0 PULSE (-10v 10v 10s 100s)

R1 a b  1
.save all @r1[i]

D1 b 0 myDiode
.model myDiode D(IS=0.1A JSW=0.2A IBV=0.3A BV=8v)

.tran 10ms 200s

.control
  run
  plot @r1[i] vs a
  plot @r1[i] vs a xlimit -250mV 0 ylimit -110mA 0
.endc

.end
