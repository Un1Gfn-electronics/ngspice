.title Working of Transistors

.model NPN0 NPN()

VC C 0 DC 0 PULSE(-1v 1v 0s 1s 1s  5s 12s)
VE E 0 DC 0 PULSE(-1v 1v 0s 1s 1s 11s 24s)
.save all @VC[i] @VE[i]

Q1 C 0 E NPN0

.control
  tran 100ms 25s
  plot C+20mV E xlimit 0ms 25s
  * plot @VC[i] @VE[i]
.endc

.end
